class coverage extends uvm_subscriber